grammar edu:umn:cs:melt:exts:ableC:checkedc;

exports edu:umn:cs:melt:exts:ableC:checkedc:concretesyntax;

exports edu:umn:cs:melt:exts:ableC:checkedc:abstractsyntax;
